`timescale 1ns / 1ps
`ifndef _param_vh_
`define _param_vh_

`define ADDR_BITS 16
`define DATA_BITS 8
`define ROM_SIZE 2048
`define MEM_SIZE (2**`ADDR_BITS)

`endif