`ifndef _opcodes_vh_
`define _opcodes_vh_

`define OP_ADD 'b00000000
`define OP_SUB 'b00000001
`define OP_MULTIPLY 'b00000010
`define OP_AND 'b00000011
`define OP_OR 'b00000100
`define OP_SROP1 'b00000101
`define OP_SLOP1 'b00000110
`define OP_NEGOP1 'b00000111
`define OP_JMP 'b00001000
`define OP_RET 'b00001001
`define OP_MVIA 'b00001011
`define OP_HALT 'b11111111

//`define OP_LDAC 'b00000001




/*`define OP_XOR 'b00000110
`define OP_OUT 'b00000111
`define OP_STAC 'b00001000
`define OP_LDA 'b00001001
`define OP_STA 'b00001010
`define OP_CMA 'b00001011
`define OP_ACA 'b00001100
*/

`endif