`ifndef _opcodes_vh_
`define _opcodes_vh_

`define OP_LDAC 'b00000001
`define OP_ADD 'b00000010
`define OP_SUB 'b00000011
`define OP_AND 'b00000100
`define OP_OR 'b00000101
`define OP_XOR 'b00000110
`define OP_OUT 'b00000111
`define OP_STAC 'b00001000
`define OP_LDA 'b00001001
`define OP_STA 'b00001010
`define OP_CMA 'b00001011
`define OP_ACA 'b00001100
`define OP_SRAC 'b00001101
`define OP_SLAC 'b00001110

`endif